
class env extends uvm_env;

endclass : env
